module fpu (a,b,fc,wf,fd,ein1,clk,clrn,ed,wd,wn,ww,st_ds,e1n,e1w, // fpu 
			e2n,e2w,e3n,e3w,e,ein2);
input clk, clrn; // clock and reset 
input [31:0] a, b; // 32-bit fp numbers 
input [4:0] fd; // fp dest reg number 
input [2:0] fc; // fp control 
input wf; // write fp regfile 
input ein1; // no_cache_stall 
input ein2; // for canceling E1 inst 
output [31:0] ed,wd; // wd: fp result 
//output [4:0] count_div,count_sqrt; // for testing 
output [4:0] e1n,e2n,e3n,wn; // reg numbers/
//output [1:0] e1c,e2c,e3c; // for testing 
output e1w,e2w,e3w,ww; // write fp regfile 
output st_ds; // stall caused by fdiv or fsqrt 
output e; // ein1 & ?st_ds 
reg [31:0] wd; 
reg [31:0] efa,efb; 
reg [4:0] e1n,e2n,e3n,wn; 
//reg [1:0] e1c,e2c,e3c; 
reg e1w0,e2w,e3w,ww,sub; 
wire [31:0] s_add;
wire [25:0] reg_x_div,reg_x_sqrt;
//wire busy_div,stall_div,busy_sqrt,stall_sqrt; 
wire fdiv = fc[2] & fc[1];
wire fsqrt = fc[2] & fc[1]; 
assign e1w = e1w0 & ein2; 
assign e = ein1;
pipelined_fadder f_add (efa,efb,sub,2'b0,s_add,clk,clrn,e); 
assign st_ds = 0;
assign ed = s_add;

always @ (negedge clrn or posedge clk) 
	if (clrn) begin // pipeline registers 
		sub <= 0; efa <= 0; efb <= 0; 
		e1w0 <= 0; e1n <= 0; 
		 e2w <= 0; e2n <= 0; 
		 e3w <= 0; e3n <= 0; 
		wd <= 0; ww <= 0; wn <= 0; 
	end else if (e) begin 
		sub <= fc[0]; efa <= a; efb <= b; 
		e1w0 <= wf; e1n <= fd; 
		 e2w <= e1w; e2n <= e1n; 
		 e3w <= e2w; e3n <= e2n; 
		wd <= ed; ww <= e3w; wn <= e3n; 
	end 
endmodule // fpu